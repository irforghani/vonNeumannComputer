Library IEEE;
Library WORK;
use STD.TEXTIO.ALL;
use IEEE.std_logic_textio.ALL;
use IEEE.STD_LOGIC_1164.ALL;
use WORK.utilities1.ALL;                                            

entity Std_Logic_Ram is 

end Std_Logic_Ram; 


architecture Behavioral of Std_Logic_Ram is 


end Behavioral; 